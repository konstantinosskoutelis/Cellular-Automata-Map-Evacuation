module weights( 
 input logic rst, 
 output logic [4095:0][12:0]weight 
); 
 always_comb begin 
weight[0] =999;
weight[1] =999;
weight[2] =999;
weight[3] =999;
weight[4] =999;
weight[5] =999;
weight[6] =999;
weight[7] =999;
weight[8] =999;
weight[9] =999;
weight[10] =999;
weight[11] =999;
weight[12] =999;
weight[13] =999;
weight[14] =999;
weight[15] =999;
weight[16] =999;
weight[17] =999;
weight[18] =999;
weight[19] =999;
weight[20] =999;
weight[21] =0;
weight[22] =999;
weight[23] =999;
weight[24] =999;
weight[25] =999;
weight[26] =999;
weight[27] =999;
weight[28] =999;
weight[29] =999;
weight[30] =999;
weight[31] =999;
weight[32] =999;
weight[33] =999;
weight[34] =999;
weight[35] =999;
weight[36] =999;
weight[37] =999;
weight[38] =999;
weight[39] =999;
weight[40] =999;
weight[41] =999;
weight[42] =999;
weight[43] =999;
weight[44] =999;
weight[45] =999;
weight[46] =999;
weight[47] =999;
weight[48] =999;
weight[49] =999;
weight[50] =999;
weight[51] =999;
weight[52] =999;
weight[53] =999;
weight[54] =999;
weight[55] =999;
weight[56] =999;
weight[57] =999;
weight[58] =999;
weight[59] =999;
weight[60] =999;
weight[61] =999;
weight[62] =999;
weight[63] =999;
weight[64] =999;
weight[65] =21;
weight[66] =20;
weight[67] =19;
weight[68] =18;
weight[69] =17;
weight[70] =16;
weight[71] =15;
weight[72] =14;
weight[73] =13;
weight[74] =12;
weight[75] =11;
weight[76] =10;
weight[77] =9;
weight[78] =8;
weight[79] =7;
weight[80] =6;
weight[81] =5;
weight[82] =4;
weight[83] =3;
weight[84] =2;
weight[85] =1;
weight[86] =2;
weight[87] =3;
weight[88] =4;
weight[89] =5;
weight[90] =6;
weight[91] =7;
weight[92] =8;
weight[93] =9;
weight[94] =10;
weight[95] =11;
weight[96] =12;
weight[97] =13;
weight[98] =14;
weight[99] =15;
weight[100] =16;
weight[101] =17;
weight[102] =18;
weight[103] =19;
weight[104] =20;
weight[105] =21;
weight[106] =22;
weight[107] =23;
weight[108] =24;
weight[109] =25;
weight[110] =26;
weight[111] =27;
weight[112] =28;
weight[113] =29;
weight[114] =30;
weight[115] =31;
weight[116] =32;
weight[117] =32;
weight[118] =31;
weight[119] =30;
weight[120] =29;
weight[121] =28;
weight[122] =27;
weight[123] =26;
weight[124] =25;
weight[125] =24;
weight[126] =23;
weight[127] =999;
weight[128] =999;
weight[129] =22;
weight[130] =21;
weight[131] =20;
weight[132] =19;
weight[133] =18;
weight[134] =17;
weight[135] =16;
weight[136] =15;
weight[137] =14;
weight[138] =13;
weight[139] =12;
weight[140] =11;
weight[141] =10;
weight[142] =9;
weight[143] =8;
weight[144] =7;
weight[145] =6;
weight[146] =5;
weight[147] =4;
weight[148] =3;
weight[149] =2;
weight[150] =3;
weight[151] =4;
weight[152] =5;
weight[153] =6;
weight[154] =7;
weight[155] =8;
weight[156] =9;
weight[157] =10;
weight[158] =11;
weight[159] =12;
weight[160] =13;
weight[161] =14;
weight[162] =15;
weight[163] =16;
weight[164] =17;
weight[165] =18;
weight[166] =19;
weight[167] =20;
weight[168] =21;
weight[169] =22;
weight[170] =23;
weight[171] =24;
weight[172] =25;
weight[173] =26;
weight[174] =27;
weight[175] =28;
weight[176] =29;
weight[177] =30;
weight[178] =31;
weight[179] =32;
weight[180] =32;
weight[181] =31;
weight[182] =30;
weight[183] =29;
weight[184] =28;
weight[185] =27;
weight[186] =26;
weight[187] =25;
weight[188] =24;
weight[189] =23;
weight[190] =22;
weight[191] =999;
weight[192] =999;
weight[193] =23;
weight[194] =22;
weight[195] =21;
weight[196] =20;
weight[197] =19;
weight[198] =18;
weight[199] =17;
weight[200] =16;
weight[201] =15;
weight[202] =14;
weight[203] =13;
weight[204] =12;
weight[205] =11;
weight[206] =10;
weight[207] =9;
weight[208] =8;
weight[209] =7;
weight[210] =6;
weight[211] =5;
weight[212] =4;
weight[213] =3;
weight[214] =4;
weight[215] =5;
weight[216] =6;
weight[217] =7;
weight[218] =8;
weight[219] =9;
weight[220] =10;
weight[221] =11;
weight[222] =12;
weight[223] =13;
weight[224] =14;
weight[225] =15;
weight[226] =16;
weight[227] =17;
weight[228] =18;
weight[229] =19;
weight[230] =20;
weight[231] =21;
weight[232] =22;
weight[233] =23;
weight[234] =24;
weight[235] =25;
weight[236] =26;
weight[237] =27;
weight[238] =28;
weight[239] =29;
weight[240] =30;
weight[241] =31;
weight[242] =32;
weight[243] =32;
weight[244] =31;
weight[245] =30;
weight[246] =29;
weight[247] =28;
weight[248] =27;
weight[249] =26;
weight[250] =25;
weight[251] =24;
weight[252] =23;
weight[253] =22;
weight[254] =21;
weight[255] =999;
weight[256] =999;
weight[257] =24;
weight[258] =23;
weight[259] =22;
weight[260] =21;
weight[261] =20;
weight[262] =19;
weight[263] =18;
weight[264] =17;
weight[265] =16;
weight[266] =15;
weight[267] =14;
weight[268] =13;
weight[269] =12;
weight[270] =11;
weight[271] =10;
weight[272] =9;
weight[273] =8;
weight[274] =7;
weight[275] =6;
weight[276] =5;
weight[277] =4;
weight[278] =5;
weight[279] =6;
weight[280] =7;
weight[281] =8;
weight[282] =9;
weight[283] =10;
weight[284] =11;
weight[285] =12;
weight[286] =13;
weight[287] =14;
weight[288] =15;
weight[289] =16;
weight[290] =17;
weight[291] =18;
weight[292] =19;
weight[293] =20;
weight[294] =21;
weight[295] =22;
weight[296] =23;
weight[297] =24;
weight[298] =25;
weight[299] =26;
weight[300] =27;
weight[301] =28;
weight[302] =29;
weight[303] =30;
weight[304] =31;
weight[305] =32;
weight[306] =32;
weight[307] =31;
weight[308] =30;
weight[309] =29;
weight[310] =28;
weight[311] =27;
weight[312] =26;
weight[313] =25;
weight[314] =24;
weight[315] =23;
weight[316] =22;
weight[317] =21;
weight[318] =20;
weight[319] =999;
weight[320] =999;
weight[321] =25;
weight[322] =24;
weight[323] =23;
weight[324] =22;
weight[325] =21;
weight[326] =20;
weight[327] =19;
weight[328] =18;
weight[329] =17;
weight[330] =16;
weight[331] =15;
weight[332] =14;
weight[333] =13;
weight[334] =12;
weight[335] =11;
weight[336] =10;
weight[337] =9;
weight[338] =8;
weight[339] =7;
weight[340] =6;
weight[341] =5;
weight[342] =6;
weight[343] =7;
weight[344] =8;
weight[345] =9;
weight[346] =10;
weight[347] =11;
weight[348] =12;
weight[349] =13;
weight[350] =14;
weight[351] =15;
weight[352] =16;
weight[353] =17;
weight[354] =18;
weight[355] =19;
weight[356] =20;
weight[357] =21;
weight[358] =22;
weight[359] =23;
weight[360] =24;
weight[361] =25;
weight[362] =26;
weight[363] =27;
weight[364] =28;
weight[365] =29;
weight[366] =30;
weight[367] =999;
weight[368] =999;
weight[369] =999;
weight[370] =999;
weight[371] =999;
weight[372] =999;
weight[373] =999;
weight[374] =999;
weight[375] =999;
weight[376] =999;
weight[377] =999;
weight[378] =999;
weight[379] =22;
weight[380] =21;
weight[381] =20;
weight[382] =19;
weight[383] =999;
weight[384] =999;
weight[385] =24;
weight[386] =25;
weight[387] =24;
weight[388] =23;
weight[389] =22;
weight[390] =21;
weight[391] =20;
weight[392] =19;
weight[393] =18;
weight[394] =17;
weight[395] =16;
weight[396] =15;
weight[397] =14;
weight[398] =13;
weight[399] =12;
weight[400] =11;
weight[401] =10;
weight[402] =9;
weight[403] =8;
weight[404] =7;
weight[405] =6;
weight[406] =7;
weight[407] =8;
weight[408] =9;
weight[409] =10;
weight[410] =11;
weight[411] =12;
weight[412] =13;
weight[413] =14;
weight[414] =15;
weight[415] =16;
weight[416] =999;
weight[417] =999;
weight[418] =19;
weight[419] =20;
weight[420] =21;
weight[421] =22;
weight[422] =23;
weight[423] =24;
weight[424] =25;
weight[425] =26;
weight[426] =27;
weight[427] =28;
weight[428] =29;
weight[429] =30;
weight[430] =31;
weight[431] =999;
weight[432] =999;
weight[433] =999;
weight[434] =999;
weight[435] =999;
weight[436] =999;
weight[437] =999;
weight[438] =999;
weight[439] =999;
weight[440] =999;
weight[441] =999;
weight[442] =999;
weight[443] =21;
weight[444] =20;
weight[445] =19;
weight[446] =18;
weight[447] =999;
weight[448] =999;
weight[449] =23;
weight[450] =24;
weight[451] =25;
weight[452] =24;
weight[453] =23;
weight[454] =22;
weight[455] =21;
weight[456] =20;
weight[457] =19;
weight[458] =18;
weight[459] =17;
weight[460] =16;
weight[461] =15;
weight[462] =14;
weight[463] =13;
weight[464] =12;
weight[465] =11;
weight[466] =10;
weight[467] =9;
weight[468] =8;
weight[469] =7;
weight[470] =8;
weight[471] =9;
weight[472] =10;
weight[473] =11;
weight[474] =12;
weight[475] =13;
weight[476] =14;
weight[477] =15;
weight[478] =16;
weight[479] =17;
weight[480] =999;
weight[481] =999;
weight[482] =20;
weight[483] =21;
weight[484] =22;
weight[485] =23;
weight[486] =24;
weight[487] =25;
weight[488] =26;
weight[489] =27;
weight[490] =28;
weight[491] =29;
weight[492] =30;
weight[493] =31;
weight[494] =32;
weight[495] =999;
weight[496] =999;
weight[497] =999;
weight[498] =999;
weight[499] =999;
weight[500] =999;
weight[501] =999;
weight[502] =999;
weight[503] =999;
weight[504] =999;
weight[505] =999;
weight[506] =999;
weight[507] =20;
weight[508] =19;
weight[509] =18;
weight[510] =17;
weight[511] =999;
weight[512] =999;
weight[513] =22;
weight[514] =23;
weight[515] =24;
weight[516] =25;
weight[517] =24;
weight[518] =23;
weight[519] =22;
weight[520] =21;
weight[521] =20;
weight[522] =19;
weight[523] =18;
weight[524] =17;
weight[525] =16;
weight[526] =15;
weight[527] =14;
weight[528] =13;
weight[529] =12;
weight[530] =11;
weight[531] =10;
weight[532] =9;
weight[533] =8;
weight[534] =9;
weight[535] =10;
weight[536] =11;
weight[537] =12;
weight[538] =13;
weight[539] =14;
weight[540] =15;
weight[541] =16;
weight[542] =17;
weight[543] =18;
weight[544] =19;
weight[545] =20;
weight[546] =21;
weight[547] =22;
weight[548] =23;
weight[549] =24;
weight[550] =25;
weight[551] =26;
weight[552] =27;
weight[553] =28;
weight[554] =29;
weight[555] =30;
weight[556] =31;
weight[557] =32;
weight[558] =32;
weight[559] =999;
weight[560] =999;
weight[561] =999;
weight[562] =999;
weight[563] =999;
weight[564] =999;
weight[565] =999;
weight[566] =999;
weight[567] =999;
weight[568] =999;
weight[569] =999;
weight[570] =999;
weight[571] =19;
weight[572] =18;
weight[573] =17;
weight[574] =16;
weight[575] =999;
weight[576] =999;
weight[577] =21;
weight[578] =22;
weight[579] =23;
weight[580] =24;
weight[581] =25;
weight[582] =24;
weight[583] =23;
weight[584] =22;
weight[585] =21;
weight[586] =20;
weight[587] =999;
weight[588] =999;
weight[589] =999;
weight[590] =16;
weight[591] =15;
weight[592] =14;
weight[593] =13;
weight[594] =12;
weight[595] =11;
weight[596] =10;
weight[597] =9;
weight[598] =10;
weight[599] =11;
weight[600] =12;
weight[601] =13;
weight[602] =14;
weight[603] =15;
weight[604] =16;
weight[605] =17;
weight[606] =18;
weight[607] =19;
weight[608] =20;
weight[609] =21;
weight[610] =22;
weight[611] =23;
weight[612] =24;
weight[613] =25;
weight[614] =26;
weight[615] =27;
weight[616] =28;
weight[617] =29;
weight[618] =30;
weight[619] =31;
weight[620] =32;
weight[621] =32;
weight[622] =31;
weight[623] =999;
weight[624] =999;
weight[625] =999;
weight[626] =999;
weight[627] =999;
weight[628] =999;
weight[629] =999;
weight[630] =999;
weight[631] =999;
weight[632] =999;
weight[633] =999;
weight[634] =999;
weight[635] =18;
weight[636] =17;
weight[637] =16;
weight[638] =15;
weight[639] =999;
weight[640] =999;
weight[641] =20;
weight[642] =21;
weight[643] =22;
weight[644] =23;
weight[645] =24;
weight[646] =25;
weight[647] =24;
weight[648] =23;
weight[649] =22;
weight[650] =21;
weight[651] =999;
weight[652] =999;
weight[653] =999;
weight[654] =17;
weight[655] =16;
weight[656] =15;
weight[657] =14;
weight[658] =13;
weight[659] =12;
weight[660] =11;
weight[661] =10;
weight[662] =11;
weight[663] =12;
weight[664] =13;
weight[665] =14;
weight[666] =15;
weight[667] =16;
weight[668] =17;
weight[669] =18;
weight[670] =19;
weight[671] =20;
weight[672] =21;
weight[673] =22;
weight[674] =23;
weight[675] =24;
weight[676] =25;
weight[677] =26;
weight[678] =27;
weight[679] =28;
weight[680] =29;
weight[681] =30;
weight[682] =31;
weight[683] =32;
weight[684] =32;
weight[685] =31;
weight[686] =30;
weight[687] =29;
weight[688] =28;
weight[689] =27;
weight[690] =26;
weight[691] =25;
weight[692] =24;
weight[693] =23;
weight[694] =22;
weight[695] =21;
weight[696] =20;
weight[697] =19;
weight[698] =18;
weight[699] =17;
weight[700] =16;
weight[701] =15;
weight[702] =14;
weight[703] =999;
weight[704] =999;
weight[705] =19;
weight[706] =20;
weight[707] =21;
weight[708] =22;
weight[709] =23;
weight[710] =24;
weight[711] =25;
weight[712] =24;
weight[713] =23;
weight[714] =22;
weight[715] =999;
weight[716] =999;
weight[717] =999;
weight[718] =18;
weight[719] =17;
weight[720] =16;
weight[721] =15;
weight[722] =14;
weight[723] =13;
weight[724] =12;
weight[725] =11;
weight[726] =12;
weight[727] =13;
weight[728] =14;
weight[729] =15;
weight[730] =16;
weight[731] =17;
weight[732] =18;
weight[733] =19;
weight[734] =20;
weight[735] =21;
weight[736] =22;
weight[737] =23;
weight[738] =24;
weight[739] =25;
weight[740] =26;
weight[741] =27;
weight[742] =28;
weight[743] =29;
weight[744] =30;
weight[745] =31;
weight[746] =32;
weight[747] =32;
weight[748] =31;
weight[749] =30;
weight[750] =29;
weight[751] =28;
weight[752] =27;
weight[753] =26;
weight[754] =25;
weight[755] =24;
weight[756] =23;
weight[757] =22;
weight[758] =21;
weight[759] =20;
weight[760] =19;
weight[761] =18;
weight[762] =17;
weight[763] =16;
weight[764] =15;
weight[765] =14;
weight[766] =13;
weight[767] =999;
weight[768] =999;
weight[769] =18;
weight[770] =19;
weight[771] =20;
weight[772] =21;
weight[773] =22;
weight[774] =23;
weight[775] =24;
weight[776] =25;
weight[777] =24;
weight[778] =23;
weight[779] =999;
weight[780] =999;
weight[781] =999;
weight[782] =19;
weight[783] =18;
weight[784] =17;
weight[785] =16;
weight[786] =15;
weight[787] =14;
weight[788] =13;
weight[789] =12;
weight[790] =13;
weight[791] =14;
weight[792] =15;
weight[793] =16;
weight[794] =17;
weight[795] =18;
weight[796] =19;
weight[797] =20;
weight[798] =21;
weight[799] =22;
weight[800] =23;
weight[801] =24;
weight[802] =25;
weight[803] =26;
weight[804] =27;
weight[805] =28;
weight[806] =29;
weight[807] =30;
weight[808] =31;
weight[809] =32;
weight[810] =32;
weight[811] =31;
weight[812] =30;
weight[813] =29;
weight[814] =28;
weight[815] =27;
weight[816] =26;
weight[817] =25;
weight[818] =24;
weight[819] =23;
weight[820] =22;
weight[821] =21;
weight[822] =20;
weight[823] =19;
weight[824] =18;
weight[825] =17;
weight[826] =16;
weight[827] =15;
weight[828] =14;
weight[829] =13;
weight[830] =12;
weight[831] =999;
weight[832] =999;
weight[833] =17;
weight[834] =18;
weight[835] =19;
weight[836] =20;
weight[837] =21;
weight[838] =22;
weight[839] =23;
weight[840] =24;
weight[841] =25;
weight[842] =24;
weight[843] =999;
weight[844] =999;
weight[845] =999;
weight[846] =20;
weight[847] =19;
weight[848] =18;
weight[849] =17;
weight[850] =16;
weight[851] =15;
weight[852] =14;
weight[853] =13;
weight[854] =14;
weight[855] =15;
weight[856] =16;
weight[857] =17;
weight[858] =18;
weight[859] =19;
weight[860] =20;
weight[861] =21;
weight[862] =22;
weight[863] =23;
weight[864] =24;
weight[865] =25;
weight[866] =26;
weight[867] =27;
weight[868] =28;
weight[869] =29;
weight[870] =30;
weight[871] =31;
weight[872] =32;
weight[873] =32;
weight[874] =31;
weight[875] =30;
weight[876] =29;
weight[877] =28;
weight[878] =27;
weight[879] =26;
weight[880] =25;
weight[881] =24;
weight[882] =23;
weight[883] =22;
weight[884] =21;
weight[885] =20;
weight[886] =19;
weight[887] =18;
weight[888] =17;
weight[889] =16;
weight[890] =15;
weight[891] =14;
weight[892] =13;
weight[893] =12;
weight[894] =11;
weight[895] =999;
weight[896] =999;
weight[897] =16;
weight[898] =17;
weight[899] =18;
weight[900] =19;
weight[901] =20;
weight[902] =21;
weight[903] =22;
weight[904] =23;
weight[905] =24;
weight[906] =25;
weight[907] =999;
weight[908] =999;
weight[909] =999;
weight[910] =21;
weight[911] =20;
weight[912] =19;
weight[913] =18;
weight[914] =17;
weight[915] =16;
weight[916] =15;
weight[917] =14;
weight[918] =15;
weight[919] =16;
weight[920] =17;
weight[921] =18;
weight[922] =19;
weight[923] =20;
weight[924] =21;
weight[925] =22;
weight[926] =23;
weight[927] =24;
weight[928] =25;
weight[929] =26;
weight[930] =27;
weight[931] =28;
weight[932] =29;
weight[933] =30;
weight[934] =31;
weight[935] =32;
weight[936] =32;
weight[937] =31;
weight[938] =30;
weight[939] =29;
weight[940] =28;
weight[941] =27;
weight[942] =26;
weight[943] =25;
weight[944] =24;
weight[945] =23;
weight[946] =22;
weight[947] =21;
weight[948] =20;
weight[949] =19;
weight[950] =18;
weight[951] =17;
weight[952] =16;
weight[953] =15;
weight[954] =14;
weight[955] =13;
weight[956] =12;
weight[957] =11;
weight[958] =10;
weight[959] =999;
weight[960] =999;
weight[961] =15;
weight[962] =16;
weight[963] =17;
weight[964] =18;
weight[965] =19;
weight[966] =20;
weight[967] =21;
weight[968] =22;
weight[969] =23;
weight[970] =24;
weight[971] =999;
weight[972] =999;
weight[973] =999;
weight[974] =22;
weight[975] =21;
weight[976] =20;
weight[977] =19;
weight[978] =18;
weight[979] =17;
weight[980] =16;
weight[981] =15;
weight[982] =16;
weight[983] =17;
weight[984] =18;
weight[985] =19;
weight[986] =20;
weight[987] =21;
weight[988] =22;
weight[989] =23;
weight[990] =24;
weight[991] =25;
weight[992] =26;
weight[993] =27;
weight[994] =28;
weight[995] =29;
weight[996] =30;
weight[997] =31;
weight[998] =32;
weight[999] =32;
weight[1000] =31;
weight[1001] =30;
weight[1002] =29;
weight[1003] =28;
weight[1004] =27;
weight[1005] =26;
weight[1006] =25;
weight[1007] =24;
weight[1008] =23;
weight[1009] =22;
weight[1010] =21;
weight[1011] =20;
weight[1012] =19;
weight[1013] =18;
weight[1014] =17;
weight[1015] =16;
weight[1016] =15;
weight[1017] =14;
weight[1018] =13;
weight[1019] =12;
weight[1020] =11;
weight[1021] =10;
weight[1022] =9;
weight[1023] =999;
weight[1024] =999;
weight[1025] =14;
weight[1026] =15;
weight[1027] =16;
weight[1028] =17;
weight[1029] =18;
weight[1030] =19;
weight[1031] =20;
weight[1032] =21;
weight[1033] =22;
weight[1034] =23;
weight[1035] =999;
weight[1036] =999;
weight[1037] =999;
weight[1038] =23;
weight[1039] =22;
weight[1040] =21;
weight[1041] =20;
weight[1042] =19;
weight[1043] =18;
weight[1044] =17;
weight[1045] =16;
weight[1046] =17;
weight[1047] =18;
weight[1048] =19;
weight[1049] =20;
weight[1050] =21;
weight[1051] =22;
weight[1052] =23;
weight[1053] =24;
weight[1054] =25;
weight[1055] =26;
weight[1056] =27;
weight[1057] =28;
weight[1058] =29;
weight[1059] =30;
weight[1060] =31;
weight[1061] =32;
weight[1062] =32;
weight[1063] =31;
weight[1064] =30;
weight[1065] =29;
weight[1066] =28;
weight[1067] =27;
weight[1068] =26;
weight[1069] =25;
weight[1070] =24;
weight[1071] =23;
weight[1072] =22;
weight[1073] =21;
weight[1074] =20;
weight[1075] =19;
weight[1076] =18;
weight[1077] =17;
weight[1078] =16;
weight[1079] =15;
weight[1080] =14;
weight[1081] =13;
weight[1082] =12;
weight[1083] =11;
weight[1084] =10;
weight[1085] =9;
weight[1086] =8;
weight[1087] =999;
weight[1088] =999;
weight[1089] =13;
weight[1090] =14;
weight[1091] =15;
weight[1092] =16;
weight[1093] =17;
weight[1094] =18;
weight[1095] =19;
weight[1096] =20;
weight[1097] =21;
weight[1098] =22;
weight[1099] =999;
weight[1100] =999;
weight[1101] =999;
weight[1102] =24;
weight[1103] =23;
weight[1104] =22;
weight[1105] =21;
weight[1106] =20;
weight[1107] =19;
weight[1108] =18;
weight[1109] =17;
weight[1110] =18;
weight[1111] =19;
weight[1112] =20;
weight[1113] =21;
weight[1114] =22;
weight[1115] =23;
weight[1116] =24;
weight[1117] =25;
weight[1118] =26;
weight[1119] =27;
weight[1120] =28;
weight[1121] =29;
weight[1122] =30;
weight[1123] =31;
weight[1124] =32;
weight[1125] =32;
weight[1126] =31;
weight[1127] =30;
weight[1128] =29;
weight[1129] =28;
weight[1130] =27;
weight[1131] =26;
weight[1132] =25;
weight[1133] =24;
weight[1134] =23;
weight[1135] =22;
weight[1136] =21;
weight[1137] =20;
weight[1138] =19;
weight[1139] =18;
weight[1140] =17;
weight[1141] =16;
weight[1142] =15;
weight[1143] =14;
weight[1144] =13;
weight[1145] =12;
weight[1146] =11;
weight[1147] =10;
weight[1148] =9;
weight[1149] =8;
weight[1150] =7;
weight[1151] =999;
weight[1152] =999;
weight[1153] =12;
weight[1154] =13;
weight[1155] =14;
weight[1156] =15;
weight[1157] =16;
weight[1158] =17;
weight[1159] =18;
weight[1160] =19;
weight[1161] =20;
weight[1162] =21;
weight[1163] =999;
weight[1164] =999;
weight[1165] =999;
weight[1166] =999;
weight[1167] =999;
weight[1168] =999;
weight[1169] =999;
weight[1170] =999;
weight[1171] =999;
weight[1172] =999;
weight[1173] =999;
weight[1174] =999;
weight[1175] =999;
weight[1176] =999;
weight[1177] =999;
weight[1178] =999;
weight[1179] =999;
weight[1180] =999;
weight[1181] =999;
weight[1182] =999;
weight[1183] =999;
weight[1184] =999;
weight[1185] =999;
weight[1186] =999;
weight[1187] =999;
weight[1188] =999;
weight[1189] =999;
weight[1190] =999;
weight[1191] =999;
weight[1192] =999;
weight[1193] =999;
weight[1194] =999;
weight[1195] =999;
weight[1196] =999;
weight[1197] =999;
weight[1198] =999;
weight[1199] =999;
weight[1200] =20;
weight[1201] =19;
weight[1202] =18;
weight[1203] =17;
weight[1204] =16;
weight[1205] =15;
weight[1206] =14;
weight[1207] =13;
weight[1208] =12;
weight[1209] =11;
weight[1210] =10;
weight[1211] =9;
weight[1212] =8;
weight[1213] =7;
weight[1214] =6;
weight[1215] =999;
weight[1216] =999;
weight[1217] =11;
weight[1218] =12;
weight[1219] =13;
weight[1220] =14;
weight[1221] =15;
weight[1222] =16;
weight[1223] =17;
weight[1224] =18;
weight[1225] =19;
weight[1226] =20;
weight[1227] =999;
weight[1228] =999;
weight[1229] =999;
weight[1230] =999;
weight[1231] =999;
weight[1232] =999;
weight[1233] =999;
weight[1234] =999;
weight[1235] =999;
weight[1236] =999;
weight[1237] =999;
weight[1238] =999;
weight[1239] =999;
weight[1240] =999;
weight[1241] =999;
weight[1242] =999;
weight[1243] =999;
weight[1244] =999;
weight[1245] =999;
weight[1246] =999;
weight[1247] =999;
weight[1248] =999;
weight[1249] =999;
weight[1250] =999;
weight[1251] =999;
weight[1252] =999;
weight[1253] =999;
weight[1254] =999;
weight[1255] =999;
weight[1256] =999;
weight[1257] =999;
weight[1258] =999;
weight[1259] =999;
weight[1260] =999;
weight[1261] =999;
weight[1262] =999;
weight[1263] =999;
weight[1264] =19;
weight[1265] =18;
weight[1266] =17;
weight[1267] =16;
weight[1268] =15;
weight[1269] =14;
weight[1270] =13;
weight[1271] =12;
weight[1272] =11;
weight[1273] =10;
weight[1274] =9;
weight[1275] =8;
weight[1276] =7;
weight[1277] =6;
weight[1278] =5;
weight[1279] =999;
weight[1280] =999;
weight[1281] =10;
weight[1282] =11;
weight[1283] =12;
weight[1284] =13;
weight[1285] =14;
weight[1286] =15;
weight[1287] =16;
weight[1288] =17;
weight[1289] =18;
weight[1290] =19;
weight[1291] =999;
weight[1292] =999;
weight[1293] =999;
weight[1294] =999;
weight[1295] =999;
weight[1296] =999;
weight[1297] =999;
weight[1298] =999;
weight[1299] =999;
weight[1300] =999;
weight[1301] =999;
weight[1302] =999;
weight[1303] =999;
weight[1304] =999;
weight[1305] =999;
weight[1306] =999;
weight[1307] =999;
weight[1308] =999;
weight[1309] =999;
weight[1310] =999;
weight[1311] =999;
weight[1312] =999;
weight[1313] =999;
weight[1314] =999;
weight[1315] =999;
weight[1316] =999;
weight[1317] =999;
weight[1318] =999;
weight[1319] =999;
weight[1320] =999;
weight[1321] =999;
weight[1322] =999;
weight[1323] =999;
weight[1324] =999;
weight[1325] =999;
weight[1326] =999;
weight[1327] =999;
weight[1328] =18;
weight[1329] =17;
weight[1330] =16;
weight[1331] =15;
weight[1332] =14;
weight[1333] =13;
weight[1334] =12;
weight[1335] =11;
weight[1336] =10;
weight[1337] =9;
weight[1338] =8;
weight[1339] =7;
weight[1340] =6;
weight[1341] =5;
weight[1342] =4;
weight[1343] =999;
weight[1344] =999;
weight[1345] =9;
weight[1346] =10;
weight[1347] =11;
weight[1348] =12;
weight[1349] =13;
weight[1350] =14;
weight[1351] =15;
weight[1352] =16;
weight[1353] =17;
weight[1354] =18;
weight[1355] =19;
weight[1356] =20;
weight[1357] =21;
weight[1358] =22;
weight[1359] =23;
weight[1360] =24;
weight[1361] =25;
weight[1362] =24;
weight[1363] =23;
weight[1364] =22;
weight[1365] =21;
weight[1366] =22;
weight[1367] =23;
weight[1368] =24;
weight[1369] =25;
weight[1370] =26;
weight[1371] =27;
weight[1372] =28;
weight[1373] =29;
weight[1374] =30;
weight[1375] =31;
weight[1376] =32;
weight[1377] =32;
weight[1378] =31;
weight[1379] =30;
weight[1380] =29;
weight[1381] =28;
weight[1382] =27;
weight[1383] =26;
weight[1384] =25;
weight[1385] =24;
weight[1386] =23;
weight[1387] =22;
weight[1388] =21;
weight[1389] =20;
weight[1390] =999;
weight[1391] =999;
weight[1392] =17;
weight[1393] =16;
weight[1394] =15;
weight[1395] =14;
weight[1396] =13;
weight[1397] =12;
weight[1398] =11;
weight[1399] =10;
weight[1400] =9;
weight[1401] =8;
weight[1402] =7;
weight[1403] =6;
weight[1404] =5;
weight[1405] =4;
weight[1406] =3;
weight[1407] =999;
weight[1408] =999;
weight[1409] =8;
weight[1410] =9;
weight[1411] =10;
weight[1412] =11;
weight[1413] =12;
weight[1414] =13;
weight[1415] =14;
weight[1416] =15;
weight[1417] =16;
weight[1418] =17;
weight[1419] =18;
weight[1420] =19;
weight[1421] =20;
weight[1422] =21;
weight[1423] =22;
weight[1424] =23;
weight[1425] =24;
weight[1426] =25;
weight[1427] =24;
weight[1428] =23;
weight[1429] =22;
weight[1430] =23;
weight[1431] =24;
weight[1432] =25;
weight[1433] =26;
weight[1434] =27;
weight[1435] =28;
weight[1436] =29;
weight[1437] =30;
weight[1438] =31;
weight[1439] =32;
weight[1440] =32;
weight[1441] =31;
weight[1442] =30;
weight[1443] =29;
weight[1444] =28;
weight[1445] =27;
weight[1446] =26;
weight[1447] =25;
weight[1448] =24;
weight[1449] =23;
weight[1450] =22;
weight[1451] =21;
weight[1452] =20;
weight[1453] =19;
weight[1454] =999;
weight[1455] =999;
weight[1456] =16;
weight[1457] =15;
weight[1458] =14;
weight[1459] =13;
weight[1460] =12;
weight[1461] =11;
weight[1462] =10;
weight[1463] =9;
weight[1464] =8;
weight[1465] =7;
weight[1466] =6;
weight[1467] =5;
weight[1468] =4;
weight[1469] =3;
weight[1470] =2;
weight[1471] =999;
weight[1472] =999;
weight[1473] =7;
weight[1474] =8;
weight[1475] =9;
weight[1476] =10;
weight[1477] =11;
weight[1478] =12;
weight[1479] =13;
weight[1480] =14;
weight[1481] =15;
weight[1482] =16;
weight[1483] =17;
weight[1484] =18;
weight[1485] =19;
weight[1486] =20;
weight[1487] =21;
weight[1488] =22;
weight[1489] =23;
weight[1490] =24;
weight[1491] =25;
weight[1492] =24;
weight[1493] =23;
weight[1494] =24;
weight[1495] =25;
weight[1496] =26;
weight[1497] =27;
weight[1498] =28;
weight[1499] =29;
weight[1500] =30;
weight[1501] =31;
weight[1502] =32;
weight[1503] =32;
weight[1504] =31;
weight[1505] =30;
weight[1506] =29;
weight[1507] =28;
weight[1508] =27;
weight[1509] =26;
weight[1510] =25;
weight[1511] =24;
weight[1512] =23;
weight[1513] =22;
weight[1514] =21;
weight[1515] =20;
weight[1516] =19;
weight[1517] =18;
weight[1518] =999;
weight[1519] =999;
weight[1520] =15;
weight[1521] =14;
weight[1522] =13;
weight[1523] =12;
weight[1524] =11;
weight[1525] =10;
weight[1526] =9;
weight[1527] =8;
weight[1528] =7;
weight[1529] =6;
weight[1530] =5;
weight[1531] =4;
weight[1532] =3;
weight[1533] =2;
weight[1534] =1;
weight[1535] =0;
weight[1536] =999;
weight[1537] =6;
weight[1538] =7;
weight[1539] =8;
weight[1540] =9;
weight[1541] =10;
weight[1542] =11;
weight[1543] =12;
weight[1544] =13;
weight[1545] =14;
weight[1546] =15;
weight[1547] =16;
weight[1548] =17;
weight[1549] =18;
weight[1550] =19;
weight[1551] =999;
weight[1552] =999;
weight[1553] =22;
weight[1554] =23;
weight[1555] =24;
weight[1556] =25;
weight[1557] =24;
weight[1558] =25;
weight[1559] =26;
weight[1560] =27;
weight[1561] =28;
weight[1562] =29;
weight[1563] =30;
weight[1564] =31;
weight[1565] =32;
weight[1566] =33;
weight[1567] =33;
weight[1568] =32;
weight[1569] =31;
weight[1570] =30;
weight[1571] =29;
weight[1572] =28;
weight[1573] =27;
weight[1574] =26;
weight[1575] =25;
weight[1576] =24;
weight[1577] =23;
weight[1578] =22;
weight[1579] =21;
weight[1580] =20;
weight[1581] =19;
weight[1582] =999;
weight[1583] =999;
weight[1584] =16;
weight[1585] =15;
weight[1586] =14;
weight[1587] =13;
weight[1588] =12;
weight[1589] =11;
weight[1590] =10;
weight[1591] =9;
weight[1592] =8;
weight[1593] =7;
weight[1594] =6;
weight[1595] =5;
weight[1596] =4;
weight[1597] =3;
weight[1598] =2;
weight[1599] =999;
weight[1600] =999;
weight[1601] =5;
weight[1602] =6;
weight[1603] =7;
weight[1604] =8;
weight[1605] =9;
weight[1606] =10;
weight[1607] =11;
weight[1608] =12;
weight[1609] =13;
weight[1610] =14;
weight[1611] =15;
weight[1612] =16;
weight[1613] =17;
weight[1614] =18;
weight[1615] =999;
weight[1616] =999;
weight[1617] =21;
weight[1618] =22;
weight[1619] =23;
weight[1620] =24;
weight[1621] =25;
weight[1622] =26;
weight[1623] =27;
weight[1624] =28;
weight[1625] =29;
weight[1626] =30;
weight[1627] =31;
weight[1628] =32;
weight[1629] =33;
weight[1630] =34;
weight[1631] =34;
weight[1632] =33;
weight[1633] =32;
weight[1634] =31;
weight[1635] =30;
weight[1636] =29;
weight[1637] =28;
weight[1638] =27;
weight[1639] =26;
weight[1640] =25;
weight[1641] =24;
weight[1642] =23;
weight[1643] =22;
weight[1644] =21;
weight[1645] =20;
weight[1646] =999;
weight[1647] =999;
weight[1648] =17;
weight[1649] =16;
weight[1650] =15;
weight[1651] =14;
weight[1652] =13;
weight[1653] =12;
weight[1654] =11;
weight[1655] =10;
weight[1656] =9;
weight[1657] =8;
weight[1658] =7;
weight[1659] =6;
weight[1660] =5;
weight[1661] =4;
weight[1662] =3;
weight[1663] =999;
weight[1664] =999;
weight[1665] =4;
weight[1666] =5;
weight[1667] =6;
weight[1668] =7;
weight[1669] =8;
weight[1670] =9;
weight[1671] =10;
weight[1672] =11;
weight[1673] =12;
weight[1674] =13;
weight[1675] =14;
weight[1676] =15;
weight[1677] =16;
weight[1678] =17;
weight[1679] =999;
weight[1680] =999;
weight[1681] =20;
weight[1682] =21;
weight[1683] =22;
weight[1684] =23;
weight[1685] =24;
weight[1686] =25;
weight[1687] =26;
weight[1688] =27;
weight[1689] =28;
weight[1690] =29;
weight[1691] =30;
weight[1692] =31;
weight[1693] =32;
weight[1694] =33;
weight[1695] =34;
weight[1696] =34;
weight[1697] =33;
weight[1698] =32;
weight[1699] =31;
weight[1700] =30;
weight[1701] =29;
weight[1702] =28;
weight[1703] =27;
weight[1704] =26;
weight[1705] =25;
weight[1706] =24;
weight[1707] =23;
weight[1708] =22;
weight[1709] =21;
weight[1710] =999;
weight[1711] =999;
weight[1712] =18;
weight[1713] =17;
weight[1714] =16;
weight[1715] =15;
weight[1716] =14;
weight[1717] =13;
weight[1718] =12;
weight[1719] =11;
weight[1720] =10;
weight[1721] =9;
weight[1722] =8;
weight[1723] =7;
weight[1724] =6;
weight[1725] =5;
weight[1726] =4;
weight[1727] =999;
weight[1728] =999;
weight[1729] =3;
weight[1730] =4;
weight[1731] =5;
weight[1732] =6;
weight[1733] =7;
weight[1734] =8;
weight[1735] =9;
weight[1736] =10;
weight[1737] =11;
weight[1738] =12;
weight[1739] =13;
weight[1740] =14;
weight[1741] =15;
weight[1742] =16;
weight[1743] =999;
weight[1744] =999;
weight[1745] =19;
weight[1746] =20;
weight[1747] =21;
weight[1748] =22;
weight[1749] =23;
weight[1750] =24;
weight[1751] =25;
weight[1752] =26;
weight[1753] =27;
weight[1754] =28;
weight[1755] =29;
weight[1756] =30;
weight[1757] =31;
weight[1758] =32;
weight[1759] =33;
weight[1760] =34;
weight[1761] =34;
weight[1762] =33;
weight[1763] =32;
weight[1764] =31;
weight[1765] =30;
weight[1766] =29;
weight[1767] =28;
weight[1768] =27;
weight[1769] =26;
weight[1770] =25;
weight[1771] =24;
weight[1772] =23;
weight[1773] =22;
weight[1774] =999;
weight[1775] =999;
weight[1776] =19;
weight[1777] =18;
weight[1778] =17;
weight[1779] =16;
weight[1780] =15;
weight[1781] =14;
weight[1782] =13;
weight[1783] =12;
weight[1784] =11;
weight[1785] =10;
weight[1786] =9;
weight[1787] =8;
weight[1788] =7;
weight[1789] =6;
weight[1790] =5;
weight[1791] =999;
weight[1792] =999;
weight[1793] =2;
weight[1794] =3;
weight[1795] =4;
weight[1796] =5;
weight[1797] =6;
weight[1798] =7;
weight[1799] =8;
weight[1800] =9;
weight[1801] =10;
weight[1802] =11;
weight[1803] =12;
weight[1804] =13;
weight[1805] =14;
weight[1806] =15;
weight[1807] =999;
weight[1808] =999;
weight[1809] =18;
weight[1810] =19;
weight[1811] =20;
weight[1812] =21;
weight[1813] =22;
weight[1814] =23;
weight[1815] =24;
weight[1816] =25;
weight[1817] =26;
weight[1818] =27;
weight[1819] =28;
weight[1820] =29;
weight[1821] =30;
weight[1822] =31;
weight[1823] =32;
weight[1824] =33;
weight[1825] =34;
weight[1826] =34;
weight[1827] =33;
weight[1828] =32;
weight[1829] =31;
weight[1830] =30;
weight[1831] =29;
weight[1832] =28;
weight[1833] =27;
weight[1834] =26;
weight[1835] =25;
weight[1836] =24;
weight[1837] =23;
weight[1838] =999;
weight[1839] =999;
weight[1840] =20;
weight[1841] =19;
weight[1842] =18;
weight[1843] =17;
weight[1844] =16;
weight[1845] =15;
weight[1846] =14;
weight[1847] =13;
weight[1848] =12;
weight[1849] =11;
weight[1850] =10;
weight[1851] =9;
weight[1852] =8;
weight[1853] =7;
weight[1854] =6;
weight[1855] =999;
weight[1856] =0;
weight[1857] =1;
weight[1858] =2;
weight[1859] =3;
weight[1860] =4;
weight[1861] =5;
weight[1862] =6;
weight[1863] =7;
weight[1864] =8;
weight[1865] =9;
weight[1866] =10;
weight[1867] =11;
weight[1868] =12;
weight[1869] =13;
weight[1870] =14;
weight[1871] =999;
weight[1872] =999;
weight[1873] =17;
weight[1874] =18;
weight[1875] =19;
weight[1876] =20;
weight[1877] =21;
weight[1878] =22;
weight[1879] =23;
weight[1880] =24;
weight[1881] =25;
weight[1882] =26;
weight[1883] =27;
weight[1884] =28;
weight[1885] =29;
weight[1886] =30;
weight[1887] =31;
weight[1888] =32;
weight[1889] =33;
weight[1890] =34;
weight[1891] =34;
weight[1892] =33;
weight[1893] =32;
weight[1894] =31;
weight[1895] =30;
weight[1896] =29;
weight[1897] =28;
weight[1898] =27;
weight[1899] =26;
weight[1900] =25;
weight[1901] =24;
weight[1902] =999;
weight[1903] =999;
weight[1904] =21;
weight[1905] =20;
weight[1906] =19;
weight[1907] =18;
weight[1908] =17;
weight[1909] =16;
weight[1910] =15;
weight[1911] =14;
weight[1912] =13;
weight[1913] =12;
weight[1914] =11;
weight[1915] =10;
weight[1916] =9;
weight[1917] =8;
weight[1918] =7;
weight[1919] =999;
weight[1920] =999;
weight[1921] =2;
weight[1922] =3;
weight[1923] =4;
weight[1924] =5;
weight[1925] =6;
weight[1926] =7;
weight[1927] =8;
weight[1928] =9;
weight[1929] =10;
weight[1930] =11;
weight[1931] =12;
weight[1932] =13;
weight[1933] =14;
weight[1934] =15;
weight[1935] =999;
weight[1936] =999;
weight[1937] =18;
weight[1938] =19;
weight[1939] =20;
weight[1940] =21;
weight[1941] =22;
weight[1942] =23;
weight[1943] =24;
weight[1944] =25;
weight[1945] =26;
weight[1946] =27;
weight[1947] =28;
weight[1948] =29;
weight[1949] =30;
weight[1950] =31;
weight[1951] =32;
weight[1952] =33;
weight[1953] =34;
weight[1954] =35;
weight[1955] =35;
weight[1956] =34;
weight[1957] =33;
weight[1958] =32;
weight[1959] =31;
weight[1960] =30;
weight[1961] =29;
weight[1962] =28;
weight[1963] =27;
weight[1964] =26;
weight[1965] =25;
weight[1966] =999;
weight[1967] =999;
weight[1968] =22;
weight[1969] =21;
weight[1970] =20;
weight[1971] =19;
weight[1972] =18;
weight[1973] =17;
weight[1974] =16;
weight[1975] =15;
weight[1976] =14;
weight[1977] =13;
weight[1978] =12;
weight[1979] =11;
weight[1980] =10;
weight[1981] =9;
weight[1982] =8;
weight[1983] =999;
weight[1984] =999;
weight[1985] =3;
weight[1986] =4;
weight[1987] =5;
weight[1988] =6;
weight[1989] =7;
weight[1990] =8;
weight[1991] =9;
weight[1992] =10;
weight[1993] =11;
weight[1994] =12;
weight[1995] =13;
weight[1996] =14;
weight[1997] =15;
weight[1998] =16;
weight[1999] =999;
weight[2000] =999;
weight[2001] =19;
weight[2002] =20;
weight[2003] =21;
weight[2004] =22;
weight[2005] =23;
weight[2006] =24;
weight[2007] =25;
weight[2008] =26;
weight[2009] =27;
weight[2010] =28;
weight[2011] =29;
weight[2012] =30;
weight[2013] =31;
weight[2014] =32;
weight[2015] =33;
weight[2016] =34;
weight[2017] =35;
weight[2018] =36;
weight[2019] =36;
weight[2020] =35;
weight[2021] =34;
weight[2022] =33;
weight[2023] =32;
weight[2024] =31;
weight[2025] =30;
weight[2026] =29;
weight[2027] =28;
weight[2028] =27;
weight[2029] =26;
weight[2030] =999;
weight[2031] =999;
weight[2032] =23;
weight[2033] =22;
weight[2034] =21;
weight[2035] =20;
weight[2036] =19;
weight[2037] =18;
weight[2038] =17;
weight[2039] =16;
weight[2040] =15;
weight[2041] =14;
weight[2042] =13;
weight[2043] =12;
weight[2044] =11;
weight[2045] =10;
weight[2046] =9;
weight[2047] =999;
weight[2048] =999;
weight[2049] =4;
weight[2050] =5;
weight[2051] =6;
weight[2052] =7;
weight[2053] =8;
weight[2054] =9;
weight[2055] =10;
weight[2056] =11;
weight[2057] =12;
weight[2058] =13;
weight[2059] =14;
weight[2060] =15;
weight[2061] =16;
weight[2062] =17;
weight[2063] =999;
weight[2064] =999;
weight[2065] =20;
weight[2066] =21;
weight[2067] =22;
weight[2068] =23;
weight[2069] =24;
weight[2070] =25;
weight[2071] =26;
weight[2072] =27;
weight[2073] =28;
weight[2074] =29;
weight[2075] =30;
weight[2076] =31;
weight[2077] =32;
weight[2078] =33;
weight[2079] =34;
weight[2080] =35;
weight[2081] =36;
weight[2082] =37;
weight[2083] =37;
weight[2084] =36;
weight[2085] =35;
weight[2086] =34;
weight[2087] =33;
weight[2088] =32;
weight[2089] =31;
weight[2090] =30;
weight[2091] =29;
weight[2092] =28;
weight[2093] =27;
weight[2094] =999;
weight[2095] =999;
weight[2096] =24;
weight[2097] =23;
weight[2098] =22;
weight[2099] =21;
weight[2100] =20;
weight[2101] =19;
weight[2102] =18;
weight[2103] =17;
weight[2104] =16;
weight[2105] =15;
weight[2106] =14;
weight[2107] =13;
weight[2108] =12;
weight[2109] =11;
weight[2110] =10;
weight[2111] =999;
weight[2112] =999;
weight[2113] =5;
weight[2114] =6;
weight[2115] =7;
weight[2116] =8;
weight[2117] =9;
weight[2118] =10;
weight[2119] =11;
weight[2120] =12;
weight[2121] =13;
weight[2122] =14;
weight[2123] =15;
weight[2124] =16;
weight[2125] =17;
weight[2126] =18;
weight[2127] =999;
weight[2128] =999;
weight[2129] =21;
weight[2130] =22;
weight[2131] =23;
weight[2132] =24;
weight[2133] =25;
weight[2134] =26;
weight[2135] =27;
weight[2136] =28;
weight[2137] =29;
weight[2138] =30;
weight[2139] =31;
weight[2140] =32;
weight[2141] =33;
weight[2142] =34;
weight[2143] =35;
weight[2144] =36;
weight[2145] =37;
weight[2146] =38;
weight[2147] =38;
weight[2148] =37;
weight[2149] =36;
weight[2150] =35;
weight[2151] =34;
weight[2152] =33;
weight[2153] =32;
weight[2154] =31;
weight[2155] =30;
weight[2156] =29;
weight[2157] =28;
weight[2158] =999;
weight[2159] =999;
weight[2160] =25;
weight[2161] =24;
weight[2162] =23;
weight[2163] =22;
weight[2164] =21;
weight[2165] =20;
weight[2166] =19;
weight[2167] =18;
weight[2168] =17;
weight[2169] =16;
weight[2170] =15;
weight[2171] =14;
weight[2172] =13;
weight[2173] =12;
weight[2174] =11;
weight[2175] =999;
weight[2176] =999;
weight[2177] =6;
weight[2178] =7;
weight[2179] =8;
weight[2180] =9;
weight[2181] =10;
weight[2182] =11;
weight[2183] =12;
weight[2184] =13;
weight[2185] =14;
weight[2186] =15;
weight[2187] =16;
weight[2188] =17;
weight[2189] =18;
weight[2190] =19;
weight[2191] =999;
weight[2192] =999;
weight[2193] =22;
weight[2194] =23;
weight[2195] =24;
weight[2196] =25;
weight[2197] =26;
weight[2198] =27;
weight[2199] =28;
weight[2200] =29;
weight[2201] =30;
weight[2202] =31;
weight[2203] =32;
weight[2204] =33;
weight[2205] =34;
weight[2206] =35;
weight[2207] =36;
weight[2208] =37;
weight[2209] =38;
weight[2210] =39;
weight[2211] =39;
weight[2212] =38;
weight[2213] =37;
weight[2214] =36;
weight[2215] =35;
weight[2216] =34;
weight[2217] =33;
weight[2218] =32;
weight[2219] =31;
weight[2220] =30;
weight[2221] =29;
weight[2222] =999;
weight[2223] =999;
weight[2224] =26;
weight[2225] =25;
weight[2226] =24;
weight[2227] =23;
weight[2228] =22;
weight[2229] =21;
weight[2230] =20;
weight[2231] =19;
weight[2232] =18;
weight[2233] =17;
weight[2234] =16;
weight[2235] =15;
weight[2236] =14;
weight[2237] =13;
weight[2238] =12;
weight[2239] =999;
weight[2240] =999;
weight[2241] =7;
weight[2242] =8;
weight[2243] =9;
weight[2244] =10;
weight[2245] =11;
weight[2246] =12;
weight[2247] =13;
weight[2248] =14;
weight[2249] =15;
weight[2250] =16;
weight[2251] =17;
weight[2252] =18;
weight[2253] =19;
weight[2254] =20;
weight[2255] =999;
weight[2256] =999;
weight[2257] =23;
weight[2258] =24;
weight[2259] =25;
weight[2260] =26;
weight[2261] =27;
weight[2262] =28;
weight[2263] =29;
weight[2264] =30;
weight[2265] =31;
weight[2266] =32;
weight[2267] =33;
weight[2268] =34;
weight[2269] =35;
weight[2270] =36;
weight[2271] =37;
weight[2272] =38;
weight[2273] =39;
weight[2274] =40;
weight[2275] =40;
weight[2276] =39;
weight[2277] =38;
weight[2278] =37;
weight[2279] =36;
weight[2280] =35;
weight[2281] =34;
weight[2282] =33;
weight[2283] =32;
weight[2284] =31;
weight[2285] =30;
weight[2286] =999;
weight[2287] =999;
weight[2288] =27;
weight[2289] =26;
weight[2290] =25;
weight[2291] =24;
weight[2292] =23;
weight[2293] =22;
weight[2294] =21;
weight[2295] =20;
weight[2296] =19;
weight[2297] =18;
weight[2298] =17;
weight[2299] =16;
weight[2300] =15;
weight[2301] =14;
weight[2302] =13;
weight[2303] =999;
weight[2304] =999;
weight[2305] =8;
weight[2306] =9;
weight[2307] =10;
weight[2308] =11;
weight[2309] =12;
weight[2310] =13;
weight[2311] =14;
weight[2312] =15;
weight[2313] =16;
weight[2314] =17;
weight[2315] =18;
weight[2316] =19;
weight[2317] =20;
weight[2318] =21;
weight[2319] =999;
weight[2320] =999;
weight[2321] =24;
weight[2322] =25;
weight[2323] =26;
weight[2324] =27;
weight[2325] =28;
weight[2326] =29;
weight[2327] =30;
weight[2328] =31;
weight[2329] =32;
weight[2330] =33;
weight[2331] =34;
weight[2332] =35;
weight[2333] =36;
weight[2334] =37;
weight[2335] =38;
weight[2336] =39;
weight[2337] =40;
weight[2338] =40;
weight[2339] =39;
weight[2340] =38;
weight[2341] =37;
weight[2342] =36;
weight[2343] =35;
weight[2344] =34;
weight[2345] =33;
weight[2346] =32;
weight[2347] =31;
weight[2348] =30;
weight[2349] =29;
weight[2350] =28;
weight[2351] =27;
weight[2352] =28;
weight[2353] =27;
weight[2354] =26;
weight[2355] =25;
weight[2356] =24;
weight[2357] =23;
weight[2358] =22;
weight[2359] =21;
weight[2360] =20;
weight[2361] =19;
weight[2362] =18;
weight[2363] =17;
weight[2364] =16;
weight[2365] =15;
weight[2366] =14;
weight[2367] =999;
weight[2368] =999;
weight[2369] =9;
weight[2370] =10;
weight[2371] =11;
weight[2372] =12;
weight[2373] =13;
weight[2374] =14;
weight[2375] =15;
weight[2376] =16;
weight[2377] =17;
weight[2378] =18;
weight[2379] =19;
weight[2380] =20;
weight[2381] =21;
weight[2382] =22;
weight[2383] =999;
weight[2384] =999;
weight[2385] =25;
weight[2386] =26;
weight[2387] =27;
weight[2388] =28;
weight[2389] =29;
weight[2390] =30;
weight[2391] =31;
weight[2392] =32;
weight[2393] =33;
weight[2394] =34;
weight[2395] =35;
weight[2396] =36;
weight[2397] =37;
weight[2398] =38;
weight[2399] =39;
weight[2400] =40;
weight[2401] =40;
weight[2402] =39;
weight[2403] =38;
weight[2404] =37;
weight[2405] =36;
weight[2406] =35;
weight[2407] =34;
weight[2408] =33;
weight[2409] =32;
weight[2410] =31;
weight[2411] =30;
weight[2412] =29;
weight[2413] =28;
weight[2414] =27;
weight[2415] =26;
weight[2416] =27;
weight[2417] =28;
weight[2418] =27;
weight[2419] =26;
weight[2420] =25;
weight[2421] =24;
weight[2422] =23;
weight[2423] =22;
weight[2424] =21;
weight[2425] =20;
weight[2426] =19;
weight[2427] =18;
weight[2428] =17;
weight[2429] =16;
weight[2430] =15;
weight[2431] =999;
weight[2432] =999;
weight[2433] =10;
weight[2434] =11;
weight[2435] =12;
weight[2436] =13;
weight[2437] =14;
weight[2438] =15;
weight[2439] =999;
weight[2440] =999;
weight[2441] =999;
weight[2442] =999;
weight[2443] =999;
weight[2444] =999;
weight[2445] =999;
weight[2446] =999;
weight[2447] =999;
weight[2448] =999;
weight[2449] =999;
weight[2450] =999;
weight[2451] =999;
weight[2452] =29;
weight[2453] =30;
weight[2454] =31;
weight[2455] =32;
weight[2456] =33;
weight[2457] =34;
weight[2458] =35;
weight[2459] =36;
weight[2460] =37;
weight[2461] =38;
weight[2462] =39;
weight[2463] =40;
weight[2464] =40;
weight[2465] =39;
weight[2466] =38;
weight[2467] =37;
weight[2468] =36;
weight[2469] =35;
weight[2470] =34;
weight[2471] =33;
weight[2472] =32;
weight[2473] =31;
weight[2474] =30;
weight[2475] =29;
weight[2476] =28;
weight[2477] =27;
weight[2478] =26;
weight[2479] =25;
weight[2480] =26;
weight[2481] =27;
weight[2482] =28;
weight[2483] =27;
weight[2484] =26;
weight[2485] =25;
weight[2486] =24;
weight[2487] =23;
weight[2488] =22;
weight[2489] =21;
weight[2490] =20;
weight[2491] =19;
weight[2492] =18;
weight[2493] =17;
weight[2494] =16;
weight[2495] =999;
weight[2496] =999;
weight[2497] =11;
weight[2498] =12;
weight[2499] =13;
weight[2500] =14;
weight[2501] =15;
weight[2502] =16;
weight[2503] =999;
weight[2504] =999;
weight[2505] =999;
weight[2506] =999;
weight[2507] =999;
weight[2508] =999;
weight[2509] =999;
weight[2510] =999;
weight[2511] =999;
weight[2512] =999;
weight[2513] =999;
weight[2514] =999;
weight[2515] =999;
weight[2516] =999;
weight[2517] =999;
weight[2518] =999;
weight[2519] =999;
weight[2520] =999;
weight[2521] =999;
weight[2522] =999;
weight[2523] =999;
weight[2524] =999;
weight[2525] =999;
weight[2526] =999;
weight[2527] =999;
weight[2528] =999;
weight[2529] =999;
weight[2530] =999;
weight[2531] =999;
weight[2532] =999;
weight[2533] =999;
weight[2534] =999;
weight[2535] =999;
weight[2536] =999;
weight[2537] =999;
weight[2538] =999;
weight[2539] =999;
weight[2540] =999;
weight[2541] =999;
weight[2542] =999;
weight[2543] =999;
weight[2544] =999;
weight[2545] =26;
weight[2546] =27;
weight[2547] =28;
weight[2548] =27;
weight[2549] =26;
weight[2550] =25;
weight[2551] =24;
weight[2552] =23;
weight[2553] =22;
weight[2554] =21;
weight[2555] =20;
weight[2556] =19;
weight[2557] =18;
weight[2558] =17;
weight[2559] =999;
weight[2560] =999;
weight[2561] =12;
weight[2562] =13;
weight[2563] =14;
weight[2564] =15;
weight[2565] =16;
weight[2566] =17;
weight[2567] =18;
weight[2568] =19;
weight[2569] =20;
weight[2570] =21;
weight[2571] =999;
weight[2572] =999;
weight[2573] =24;
weight[2574] =25;
weight[2575] =26;
weight[2576] =27;
weight[2577] =28;
weight[2578] =29;
weight[2579] =30;
weight[2580] =31;
weight[2581] =32;
weight[2582] =33;
weight[2583] =34;
weight[2584] =35;
weight[2585] =36;
weight[2586] =37;
weight[2587] =38;
weight[2588] =39;
weight[2589] =40;
weight[2590] =40;
weight[2591] =39;
weight[2592] =38;
weight[2593] =37;
weight[2594] =36;
weight[2595] =999;
weight[2596] =999;
weight[2597] =999;
weight[2598] =999;
weight[2599] =999;
weight[2600] =999;
weight[2601] =999;
weight[2602] =999;
weight[2603] =999;
weight[2604] =999;
weight[2605] =999;
weight[2606] =999;
weight[2607] =999;
weight[2608] =999;
weight[2609] =25;
weight[2610] =26;
weight[2611] =27;
weight[2612] =28;
weight[2613] =27;
weight[2614] =26;
weight[2615] =25;
weight[2616] =24;
weight[2617] =23;
weight[2618] =22;
weight[2619] =21;
weight[2620] =20;
weight[2621] =19;
weight[2622] =18;
weight[2623] =999;
weight[2624] =999;
weight[2625] =13;
weight[2626] =14;
weight[2627] =15;
weight[2628] =16;
weight[2629] =17;
weight[2630] =18;
weight[2631] =19;
weight[2632] =20;
weight[2633] =21;
weight[2634] =22;
weight[2635] =999;
weight[2636] =999;
weight[2637] =25;
weight[2638] =26;
weight[2639] =27;
weight[2640] =28;
weight[2641] =29;
weight[2642] =30;
weight[2643] =31;
weight[2644] =32;
weight[2645] =33;
weight[2646] =34;
weight[2647] =35;
weight[2648] =36;
weight[2649] =37;
weight[2650] =38;
weight[2651] =39;
weight[2652] =40;
weight[2653] =40;
weight[2654] =39;
weight[2655] =38;
weight[2656] =37;
weight[2657] =36;
weight[2658] =35;
weight[2659] =999;
weight[2660] =999;
weight[2661] =999;
weight[2662] =999;
weight[2663] =999;
weight[2664] =999;
weight[2665] =999;
weight[2666] =999;
weight[2667] =999;
weight[2668] =999;
weight[2669] =999;
weight[2670] =999;
weight[2671] =999;
weight[2672] =999;
weight[2673] =24;
weight[2674] =25;
weight[2675] =26;
weight[2676] =27;
weight[2677] =28;
weight[2678] =27;
weight[2679] =26;
weight[2680] =25;
weight[2681] =24;
weight[2682] =23;
weight[2683] =22;
weight[2684] =21;
weight[2685] =20;
weight[2686] =19;
weight[2687] =999;
weight[2688] =999;
weight[2689] =14;
weight[2690] =15;
weight[2691] =16;
weight[2692] =17;
weight[2693] =18;
weight[2694] =19;
weight[2695] =20;
weight[2696] =21;
weight[2697] =22;
weight[2698] =23;
weight[2699] =999;
weight[2700] =999;
weight[2701] =26;
weight[2702] =27;
weight[2703] =28;
weight[2704] =29;
weight[2705] =30;
weight[2706] =31;
weight[2707] =32;
weight[2708] =33;
weight[2709] =34;
weight[2710] =35;
weight[2711] =36;
weight[2712] =37;
weight[2713] =38;
weight[2714] =39;
weight[2715] =40;
weight[2716] =40;
weight[2717] =39;
weight[2718] =38;
weight[2719] =37;
weight[2720] =36;
weight[2721] =35;
weight[2722] =34;
weight[2723] =999;
weight[2724] =999;
weight[2725] =999;
weight[2726] =999;
weight[2727] =999;
weight[2728] =999;
weight[2729] =999;
weight[2730] =999;
weight[2731] =999;
weight[2732] =999;
weight[2733] =999;
weight[2734] =999;
weight[2735] =999;
weight[2736] =999;
weight[2737] =23;
weight[2738] =24;
weight[2739] =25;
weight[2740] =26;
weight[2741] =27;
weight[2742] =28;
weight[2743] =27;
weight[2744] =26;
weight[2745] =25;
weight[2746] =24;
weight[2747] =23;
weight[2748] =22;
weight[2749] =21;
weight[2750] =20;
weight[2751] =999;
weight[2752] =999;
weight[2753] =15;
weight[2754] =16;
weight[2755] =17;
weight[2756] =18;
weight[2757] =19;
weight[2758] =20;
weight[2759] =21;
weight[2760] =22;
weight[2761] =23;
weight[2762] =24;
weight[2763] =999;
weight[2764] =999;
weight[2765] =27;
weight[2766] =28;
weight[2767] =29;
weight[2768] =30;
weight[2769] =31;
weight[2770] =32;
weight[2771] =33;
weight[2772] =34;
weight[2773] =35;
weight[2774] =36;
weight[2775] =37;
weight[2776] =38;
weight[2777] =39;
weight[2778] =40;
weight[2779] =40;
weight[2780] =39;
weight[2781] =38;
weight[2782] =37;
weight[2783] =36;
weight[2784] =35;
weight[2785] =34;
weight[2786] =33;
weight[2787] =999;
weight[2788] =999;
weight[2789] =999;
weight[2790] =999;
weight[2791] =999;
weight[2792] =999;
weight[2793] =999;
weight[2794] =999;
weight[2795] =999;
weight[2796] =999;
weight[2797] =999;
weight[2798] =999;
weight[2799] =999;
weight[2800] =999;
weight[2801] =22;
weight[2802] =23;
weight[2803] =24;
weight[2804] =25;
weight[2805] =26;
weight[2806] =27;
weight[2807] =28;
weight[2808] =27;
weight[2809] =26;
weight[2810] =25;
weight[2811] =24;
weight[2812] =23;
weight[2813] =22;
weight[2814] =21;
weight[2815] =999;
weight[2816] =999;
weight[2817] =16;
weight[2818] =17;
weight[2819] =18;
weight[2820] =19;
weight[2821] =20;
weight[2822] =21;
weight[2823] =22;
weight[2824] =23;
weight[2825] =24;
weight[2826] =25;
weight[2827] =999;
weight[2828] =999;
weight[2829] =28;
weight[2830] =29;
weight[2831] =30;
weight[2832] =31;
weight[2833] =32;
weight[2834] =33;
weight[2835] =34;
weight[2836] =35;
weight[2837] =36;
weight[2838] =37;
weight[2839] =38;
weight[2840] =39;
weight[2841] =40;
weight[2842] =40;
weight[2843] =39;
weight[2844] =38;
weight[2845] =37;
weight[2846] =36;
weight[2847] =35;
weight[2848] =34;
weight[2849] =33;
weight[2850] =32;
weight[2851] =999;
weight[2852] =999;
weight[2853] =999;
weight[2854] =999;
weight[2855] =999;
weight[2856] =999;
weight[2857] =999;
weight[2858] =999;
weight[2859] =999;
weight[2860] =999;
weight[2861] =999;
weight[2862] =999;
weight[2863] =999;
weight[2864] =999;
weight[2865] =21;
weight[2866] =22;
weight[2867] =23;
weight[2868] =24;
weight[2869] =25;
weight[2870] =26;
weight[2871] =27;
weight[2872] =28;
weight[2873] =27;
weight[2874] =26;
weight[2875] =25;
weight[2876] =24;
weight[2877] =23;
weight[2878] =22;
weight[2879] =999;
weight[2880] =999;
weight[2881] =17;
weight[2882] =18;
weight[2883] =19;
weight[2884] =20;
weight[2885] =21;
weight[2886] =22;
weight[2887] =23;
weight[2888] =24;
weight[2889] =25;
weight[2890] =26;
weight[2891] =999;
weight[2892] =999;
weight[2893] =29;
weight[2894] =30;
weight[2895] =31;
weight[2896] =32;
weight[2897] =33;
weight[2898] =34;
weight[2899] =35;
weight[2900] =36;
weight[2901] =37;
weight[2902] =38;
weight[2903] =39;
weight[2904] =40;
weight[2905] =40;
weight[2906] =39;
weight[2907] =38;
weight[2908] =37;
weight[2909] =36;
weight[2910] =35;
weight[2911] =34;
weight[2912] =33;
weight[2913] =32;
weight[2914] =31;
weight[2915] =999;
weight[2916] =999;
weight[2917] =999;
weight[2918] =999;
weight[2919] =999;
weight[2920] =999;
weight[2921] =999;
weight[2922] =999;
weight[2923] =999;
weight[2924] =999;
weight[2925] =999;
weight[2926] =999;
weight[2927] =999;
weight[2928] =999;
weight[2929] =20;
weight[2930] =21;
weight[2931] =22;
weight[2932] =23;
weight[2933] =24;
weight[2934] =25;
weight[2935] =26;
weight[2936] =27;
weight[2937] =28;
weight[2938] =27;
weight[2939] =26;
weight[2940] =25;
weight[2941] =24;
weight[2942] =23;
weight[2943] =999;
weight[2944] =999;
weight[2945] =18;
weight[2946] =19;
weight[2947] =20;
weight[2948] =21;
weight[2949] =22;
weight[2950] =23;
weight[2951] =24;
weight[2952] =25;
weight[2953] =26;
weight[2954] =27;
weight[2955] =999;
weight[2956] =999;
weight[2957] =30;
weight[2958] =31;
weight[2959] =32;
weight[2960] =33;
weight[2961] =34;
weight[2962] =35;
weight[2963] =36;
weight[2964] =37;
weight[2965] =38;
weight[2966] =39;
weight[2967] =40;
weight[2968] =40;
weight[2969] =39;
weight[2970] =38;
weight[2971] =37;
weight[2972] =36;
weight[2973] =35;
weight[2974] =34;
weight[2975] =33;
weight[2976] =32;
weight[2977] =31;
weight[2978] =30;
weight[2979] =999;
weight[2980] =999;
weight[2981] =999;
weight[2982] =999;
weight[2983] =999;
weight[2984] =999;
weight[2985] =999;
weight[2986] =999;
weight[2987] =999;
weight[2988] =999;
weight[2989] =999;
weight[2990] =999;
weight[2991] =999;
weight[2992] =999;
weight[2993] =19;
weight[2994] =20;
weight[2995] =21;
weight[2996] =22;
weight[2997] =23;
weight[2998] =24;
weight[2999] =25;
weight[3000] =26;
weight[3001] =27;
weight[3002] =28;
weight[3003] =27;
weight[3004] =26;
weight[3005] =25;
weight[3006] =24;
weight[3007] =999;
weight[3008] =999;
weight[3009] =19;
weight[3010] =20;
weight[3011] =21;
weight[3012] =22;
weight[3013] =23;
weight[3014] =24;
weight[3015] =25;
weight[3016] =26;
weight[3017] =27;
weight[3018] =28;
weight[3019] =999;
weight[3020] =999;
weight[3021] =31;
weight[3022] =32;
weight[3023] =33;
weight[3024] =34;
weight[3025] =35;
weight[3026] =36;
weight[3027] =37;
weight[3028] =38;
weight[3029] =39;
weight[3030] =40;
weight[3031] =40;
weight[3032] =39;
weight[3033] =38;
weight[3034] =37;
weight[3035] =36;
weight[3036] =35;
weight[3037] =34;
weight[3038] =33;
weight[3039] =32;
weight[3040] =31;
weight[3041] =30;
weight[3042] =29;
weight[3043] =999;
weight[3044] =999;
weight[3045] =999;
weight[3046] =999;
weight[3047] =999;
weight[3048] =999;
weight[3049] =999;
weight[3050] =999;
weight[3051] =999;
weight[3052] =999;
weight[3053] =999;
weight[3054] =999;
weight[3055] =999;
weight[3056] =999;
weight[3057] =18;
weight[3058] =19;
weight[3059] =20;
weight[3060] =21;
weight[3061] =22;
weight[3062] =23;
weight[3063] =24;
weight[3064] =25;
weight[3065] =26;
weight[3066] =27;
weight[3067] =28;
weight[3068] =27;
weight[3069] =26;
weight[3070] =25;
weight[3071] =999;
weight[3072] =999;
weight[3073] =20;
weight[3074] =21;
weight[3075] =22;
weight[3076] =23;
weight[3077] =24;
weight[3078] =25;
weight[3079] =26;
weight[3080] =27;
weight[3081] =28;
weight[3082] =29;
weight[3083] =999;
weight[3084] =999;
weight[3085] =32;
weight[3086] =33;
weight[3087] =34;
weight[3088] =35;
weight[3089] =36;
weight[3090] =37;
weight[3091] =38;
weight[3092] =39;
weight[3093] =40;
weight[3094] =40;
weight[3095] =39;
weight[3096] =38;
weight[3097] =37;
weight[3098] =36;
weight[3099] =35;
weight[3100] =34;
weight[3101] =33;
weight[3102] =32;
weight[3103] =31;
weight[3104] =30;
weight[3105] =29;
weight[3106] =28;
weight[3107] =999;
weight[3108] =999;
weight[3109] =999;
weight[3110] =999;
weight[3111] =999;
weight[3112] =999;
weight[3113] =999;
weight[3114] =999;
weight[3115] =999;
weight[3116] =999;
weight[3117] =999;
weight[3118] =999;
weight[3119] =999;
weight[3120] =999;
weight[3121] =17;
weight[3122] =18;
weight[3123] =19;
weight[3124] =20;
weight[3125] =21;
weight[3126] =22;
weight[3127] =23;
weight[3128] =24;
weight[3129] =25;
weight[3130] =26;
weight[3131] =27;
weight[3132] =28;
weight[3133] =27;
weight[3134] =26;
weight[3135] =999;
weight[3136] =999;
weight[3137] =21;
weight[3138] =22;
weight[3139] =23;
weight[3140] =24;
weight[3141] =25;
weight[3142] =26;
weight[3143] =27;
weight[3144] =28;
weight[3145] =29;
weight[3146] =30;
weight[3147] =999;
weight[3148] =999;
weight[3149] =33;
weight[3150] =34;
weight[3151] =35;
weight[3152] =36;
weight[3153] =37;
weight[3154] =38;
weight[3155] =39;
weight[3156] =40;
weight[3157] =40;
weight[3158] =39;
weight[3159] =38;
weight[3160] =37;
weight[3161] =36;
weight[3162] =35;
weight[3163] =34;
weight[3164] =33;
weight[3165] =32;
weight[3166] =31;
weight[3167] =30;
weight[3168] =29;
weight[3169] =28;
weight[3170] =27;
weight[3171] =999;
weight[3172] =999;
weight[3173] =999;
weight[3174] =999;
weight[3175] =999;
weight[3176] =999;
weight[3177] =999;
weight[3178] =999;
weight[3179] =999;
weight[3180] =999;
weight[3181] =999;
weight[3182] =999;
weight[3183] =999;
weight[3184] =999;
weight[3185] =16;
weight[3186] =17;
weight[3187] =18;
weight[3188] =19;
weight[3189] =20;
weight[3190] =21;
weight[3191] =22;
weight[3192] =23;
weight[3193] =24;
weight[3194] =25;
weight[3195] =26;
weight[3196] =27;
weight[3197] =28;
weight[3198] =27;
weight[3199] =999;
weight[3200] =999;
weight[3201] =22;
weight[3202] =23;
weight[3203] =24;
weight[3204] =25;
weight[3205] =26;
weight[3206] =27;
weight[3207] =28;
weight[3208] =29;
weight[3209] =30;
weight[3210] =31;
weight[3211] =999;
weight[3212] =999;
weight[3213] =34;
weight[3214] =35;
weight[3215] =36;
weight[3216] =37;
weight[3217] =38;
weight[3218] =39;
weight[3219] =40;
weight[3220] =40;
weight[3221] =39;
weight[3222] =38;
weight[3223] =37;
weight[3224] =36;
weight[3225] =35;
weight[3226] =34;
weight[3227] =33;
weight[3228] =32;
weight[3229] =31;
weight[3230] =30;
weight[3231] =29;
weight[3232] =28;
weight[3233] =27;
weight[3234] =26;
weight[3235] =999;
weight[3236] =999;
weight[3237] =999;
weight[3238] =999;
weight[3239] =999;
weight[3240] =999;
weight[3241] =999;
weight[3242] =999;
weight[3243] =999;
weight[3244] =999;
weight[3245] =999;
weight[3246] =999;
weight[3247] =999;
weight[3248] =999;
weight[3249] =15;
weight[3250] =16;
weight[3251] =17;
weight[3252] =18;
weight[3253] =19;
weight[3254] =20;
weight[3255] =21;
weight[3256] =22;
weight[3257] =23;
weight[3258] =24;
weight[3259] =25;
weight[3260] =26;
weight[3261] =27;
weight[3262] =28;
weight[3263] =999;
weight[3264] =999;
weight[3265] =23;
weight[3266] =24;
weight[3267] =25;
weight[3268] =26;
weight[3269] =27;
weight[3270] =28;
weight[3271] =29;
weight[3272] =30;
weight[3273] =31;
weight[3274] =32;
weight[3275] =999;
weight[3276] =999;
weight[3277] =35;
weight[3278] =36;
weight[3279] =37;
weight[3280] =38;
weight[3281] =39;
weight[3282] =40;
weight[3283] =40;
weight[3284] =39;
weight[3285] =38;
weight[3286] =37;
weight[3287] =36;
weight[3288] =35;
weight[3289] =34;
weight[3290] =33;
weight[3291] =32;
weight[3292] =31;
weight[3293] =30;
weight[3294] =29;
weight[3295] =28;
weight[3296] =27;
weight[3297] =26;
weight[3298] =25;
weight[3299] =999;
weight[3300] =999;
weight[3301] =999;
weight[3302] =999;
weight[3303] =999;
weight[3304] =999;
weight[3305] =999;
weight[3306] =999;
weight[3307] =999;
weight[3308] =999;
weight[3309] =999;
weight[3310] =999;
weight[3311] =999;
weight[3312] =999;
weight[3313] =14;
weight[3314] =15;
weight[3315] =16;
weight[3316] =17;
weight[3317] =18;
weight[3318] =19;
weight[3319] =20;
weight[3320] =21;
weight[3321] =22;
weight[3322] =23;
weight[3323] =24;
weight[3324] =25;
weight[3325] =26;
weight[3326] =27;
weight[3327] =999;
weight[3328] =999;
weight[3329] =24;
weight[3330] =25;
weight[3331] =26;
weight[3332] =27;
weight[3333] =28;
weight[3334] =29;
weight[3335] =30;
weight[3336] =31;
weight[3337] =32;
weight[3338] =33;
weight[3339] =999;
weight[3340] =999;
weight[3341] =36;
weight[3342] =37;
weight[3343] =38;
weight[3344] =39;
weight[3345] =40;
weight[3346] =40;
weight[3347] =39;
weight[3348] =38;
weight[3349] =37;
weight[3350] =36;
weight[3351] =35;
weight[3352] =34;
weight[3353] =33;
weight[3354] =32;
weight[3355] =31;
weight[3356] =30;
weight[3357] =29;
weight[3358] =28;
weight[3359] =27;
weight[3360] =26;
weight[3361] =25;
weight[3362] =24;
weight[3363] =999;
weight[3364] =999;
weight[3365] =999;
weight[3366] =999;
weight[3367] =999;
weight[3368] =999;
weight[3369] =999;
weight[3370] =999;
weight[3371] =999;
weight[3372] =999;
weight[3373] =999;
weight[3374] =999;
weight[3375] =999;
weight[3376] =999;
weight[3377] =13;
weight[3378] =14;
weight[3379] =15;
weight[3380] =16;
weight[3381] =17;
weight[3382] =18;
weight[3383] =19;
weight[3384] =20;
weight[3385] =21;
weight[3386] =22;
weight[3387] =23;
weight[3388] =24;
weight[3389] =25;
weight[3390] =26;
weight[3391] =999;
weight[3392] =999;
weight[3393] =25;
weight[3394] =26;
weight[3395] =27;
weight[3396] =28;
weight[3397] =29;
weight[3398] =30;
weight[3399] =31;
weight[3400] =32;
weight[3401] =33;
weight[3402] =34;
weight[3403] =999;
weight[3404] =999;
weight[3405] =37;
weight[3406] =38;
weight[3407] =39;
weight[3408] =40;
weight[3409] =40;
weight[3410] =39;
weight[3411] =38;
weight[3412] =37;
weight[3413] =36;
weight[3414] =35;
weight[3415] =34;
weight[3416] =33;
weight[3417] =32;
weight[3418] =31;
weight[3419] =30;
weight[3420] =29;
weight[3421] =28;
weight[3422] =27;
weight[3423] =26;
weight[3424] =25;
weight[3425] =24;
weight[3426] =23;
weight[3427] =999;
weight[3428] =999;
weight[3429] =999;
weight[3430] =999;
weight[3431] =999;
weight[3432] =999;
weight[3433] =999;
weight[3434] =999;
weight[3435] =999;
weight[3436] =999;
weight[3437] =999;
weight[3438] =999;
weight[3439] =999;
weight[3440] =999;
weight[3441] =12;
weight[3442] =13;
weight[3443] =14;
weight[3444] =15;
weight[3445] =16;
weight[3446] =17;
weight[3447] =18;
weight[3448] =19;
weight[3449] =20;
weight[3450] =21;
weight[3451] =22;
weight[3452] =23;
weight[3453] =24;
weight[3454] =25;
weight[3455] =999;
weight[3456] =999;
weight[3457] =26;
weight[3458] =27;
weight[3459] =28;
weight[3460] =29;
weight[3461] =30;
weight[3462] =31;
weight[3463] =32;
weight[3464] =33;
weight[3465] =34;
weight[3466] =35;
weight[3467] =999;
weight[3468] =999;
weight[3469] =38;
weight[3470] =39;
weight[3471] =40;
weight[3472] =40;
weight[3473] =39;
weight[3474] =38;
weight[3475] =37;
weight[3476] =36;
weight[3477] =35;
weight[3478] =34;
weight[3479] =33;
weight[3480] =32;
weight[3481] =31;
weight[3482] =30;
weight[3483] =29;
weight[3484] =28;
weight[3485] =27;
weight[3486] =26;
weight[3487] =25;
weight[3488] =24;
weight[3489] =23;
weight[3490] =22;
weight[3491] =21;
weight[3492] =20;
weight[3493] =19;
weight[3494] =18;
weight[3495] =17;
weight[3496] =16;
weight[3497] =15;
weight[3498] =14;
weight[3499] =13;
weight[3500] =12;
weight[3501] =11;
weight[3502] =10;
weight[3503] =9;
weight[3504] =10;
weight[3505] =11;
weight[3506] =12;
weight[3507] =13;
weight[3508] =14;
weight[3509] =15;
weight[3510] =16;
weight[3511] =17;
weight[3512] =18;
weight[3513] =19;
weight[3514] =20;
weight[3515] =21;
weight[3516] =22;
weight[3517] =23;
weight[3518] =24;
weight[3519] =999;
weight[3520] =999;
weight[3521] =27;
weight[3522] =28;
weight[3523] =29;
weight[3524] =30;
weight[3525] =31;
weight[3526] =32;
weight[3527] =33;
weight[3528] =34;
weight[3529] =35;
weight[3530] =36;
weight[3531] =37;
weight[3532] =38;
weight[3533] =39;
weight[3534] =40;
weight[3535] =40;
weight[3536] =39;
weight[3537] =38;
weight[3538] =37;
weight[3539] =36;
weight[3540] =35;
weight[3541] =34;
weight[3542] =33;
weight[3543] =32;
weight[3544] =31;
weight[3545] =30;
weight[3546] =29;
weight[3547] =28;
weight[3548] =27;
weight[3549] =26;
weight[3550] =25;
weight[3551] =24;
weight[3552] =23;
weight[3553] =22;
weight[3554] =21;
weight[3555] =20;
weight[3556] =19;
weight[3557] =18;
weight[3558] =17;
weight[3559] =16;
weight[3560] =15;
weight[3561] =14;
weight[3562] =13;
weight[3563] =12;
weight[3564] =11;
weight[3565] =10;
weight[3566] =9;
weight[3567] =8;
weight[3568] =9;
weight[3569] =10;
weight[3570] =11;
weight[3571] =12;
weight[3572] =13;
weight[3573] =14;
weight[3574] =15;
weight[3575] =16;
weight[3576] =17;
weight[3577] =18;
weight[3578] =19;
weight[3579] =20;
weight[3580] =21;
weight[3581] =22;
weight[3582] =23;
weight[3583] =999;
weight[3584] =999;
weight[3585] =28;
weight[3586] =29;
weight[3587] =30;
weight[3588] =31;
weight[3589] =32;
weight[3590] =33;
weight[3591] =34;
weight[3592] =35;
weight[3593] =36;
weight[3594] =37;
weight[3595] =38;
weight[3596] =39;
weight[3597] =40;
weight[3598] =40;
weight[3599] =39;
weight[3600] =38;
weight[3601] =37;
weight[3602] =36;
weight[3603] =35;
weight[3604] =34;
weight[3605] =33;
weight[3606] =32;
weight[3607] =31;
weight[3608] =30;
weight[3609] =29;
weight[3610] =28;
weight[3611] =27;
weight[3612] =26;
weight[3613] =25;
weight[3614] =24;
weight[3615] =23;
weight[3616] =22;
weight[3617] =21;
weight[3618] =20;
weight[3619] =19;
weight[3620] =18;
weight[3621] =17;
weight[3622] =16;
weight[3623] =15;
weight[3624] =14;
weight[3625] =13;
weight[3626] =12;
weight[3627] =11;
weight[3628] =10;
weight[3629] =9;
weight[3630] =8;
weight[3631] =7;
weight[3632] =8;
weight[3633] =9;
weight[3634] =10;
weight[3635] =11;
weight[3636] =12;
weight[3637] =13;
weight[3638] =14;
weight[3639] =15;
weight[3640] =16;
weight[3641] =17;
weight[3642] =18;
weight[3643] =19;
weight[3644] =20;
weight[3645] =21;
weight[3646] =22;
weight[3647] =999;
weight[3648] =999;
weight[3649] =29;
weight[3650] =30;
weight[3651] =31;
weight[3652] =32;
weight[3653] =33;
weight[3654] =34;
weight[3655] =35;
weight[3656] =36;
weight[3657] =37;
weight[3658] =38;
weight[3659] =39;
weight[3660] =40;
weight[3661] =40;
weight[3662] =39;
weight[3663] =38;
weight[3664] =37;
weight[3665] =36;
weight[3666] =35;
weight[3667] =34;
weight[3668] =33;
weight[3669] =32;
weight[3670] =31;
weight[3671] =30;
weight[3672] =29;
weight[3673] =28;
weight[3674] =27;
weight[3675] =26;
weight[3676] =25;
weight[3677] =24;
weight[3678] =23;
weight[3679] =22;
weight[3680] =21;
weight[3681] =20;
weight[3682] =19;
weight[3683] =18;
weight[3684] =17;
weight[3685] =16;
weight[3686] =15;
weight[3687] =14;
weight[3688] =13;
weight[3689] =12;
weight[3690] =11;
weight[3691] =10;
weight[3692] =9;
weight[3693] =8;
weight[3694] =7;
weight[3695] =6;
weight[3696] =7;
weight[3697] =8;
weight[3698] =9;
weight[3699] =10;
weight[3700] =11;
weight[3701] =12;
weight[3702] =13;
weight[3703] =14;
weight[3704] =15;
weight[3705] =16;
weight[3706] =17;
weight[3707] =18;
weight[3708] =19;
weight[3709] =20;
weight[3710] =21;
weight[3711] =999;
weight[3712] =999;
weight[3713] =30;
weight[3714] =31;
weight[3715] =32;
weight[3716] =33;
weight[3717] =34;
weight[3718] =35;
weight[3719] =36;
weight[3720] =37;
weight[3721] =38;
weight[3722] =39;
weight[3723] =40;
weight[3724] =40;
weight[3725] =39;
weight[3726] =38;
weight[3727] =37;
weight[3728] =36;
weight[3729] =35;
weight[3730] =34;
weight[3731] =33;
weight[3732] =32;
weight[3733] =31;
weight[3734] =30;
weight[3735] =29;
weight[3736] =28;
weight[3737] =27;
weight[3738] =26;
weight[3739] =25;
weight[3740] =24;
weight[3741] =23;
weight[3742] =22;
weight[3743] =21;
weight[3744] =20;
weight[3745] =19;
weight[3746] =18;
weight[3747] =17;
weight[3748] =16;
weight[3749] =15;
weight[3750] =14;
weight[3751] =13;
weight[3752] =12;
weight[3753] =11;
weight[3754] =10;
weight[3755] =9;
weight[3756] =8;
weight[3757] =7;
weight[3758] =6;
weight[3759] =5;
weight[3760] =6;
weight[3761] =7;
weight[3762] =8;
weight[3763] =9;
weight[3764] =10;
weight[3765] =11;
weight[3766] =12;
weight[3767] =13;
weight[3768] =14;
weight[3769] =15;
weight[3770] =16;
weight[3771] =17;
weight[3772] =18;
weight[3773] =19;
weight[3774] =20;
weight[3775] =999;
weight[3776] =999;
weight[3777] =31;
weight[3778] =32;
weight[3779] =33;
weight[3780] =34;
weight[3781] =35;
weight[3782] =36;
weight[3783] =37;
weight[3784] =38;
weight[3785] =39;
weight[3786] =40;
weight[3787] =40;
weight[3788] =39;
weight[3789] =38;
weight[3790] =37;
weight[3791] =36;
weight[3792] =35;
weight[3793] =34;
weight[3794] =33;
weight[3795] =32;
weight[3796] =31;
weight[3797] =30;
weight[3798] =29;
weight[3799] =28;
weight[3800] =27;
weight[3801] =26;
weight[3802] =25;
weight[3803] =24;
weight[3804] =23;
weight[3805] =22;
weight[3806] =21;
weight[3807] =20;
weight[3808] =19;
weight[3809] =18;
weight[3810] =17;
weight[3811] =16;
weight[3812] =15;
weight[3813] =14;
weight[3814] =13;
weight[3815] =12;
weight[3816] =11;
weight[3817] =10;
weight[3818] =9;
weight[3819] =8;
weight[3820] =7;
weight[3821] =6;
weight[3822] =5;
weight[3823] =4;
weight[3824] =5;
weight[3825] =6;
weight[3826] =7;
weight[3827] =8;
weight[3828] =9;
weight[3829] =10;
weight[3830] =11;
weight[3831] =12;
weight[3832] =13;
weight[3833] =14;
weight[3834] =15;
weight[3835] =16;
weight[3836] =17;
weight[3837] =18;
weight[3838] =19;
weight[3839] =999;
weight[3840] =999;
weight[3841] =32;
weight[3842] =33;
weight[3843] =34;
weight[3844] =35;
weight[3845] =36;
weight[3846] =37;
weight[3847] =38;
weight[3848] =39;
weight[3849] =40;
weight[3850] =40;
weight[3851] =39;
weight[3852] =38;
weight[3853] =37;
weight[3854] =36;
weight[3855] =35;
weight[3856] =34;
weight[3857] =33;
weight[3858] =32;
weight[3859] =31;
weight[3860] =30;
weight[3861] =29;
weight[3862] =28;
weight[3863] =27;
weight[3864] =26;
weight[3865] =25;
weight[3866] =24;
weight[3867] =23;
weight[3868] =22;
weight[3869] =21;
weight[3870] =20;
weight[3871] =19;
weight[3872] =18;
weight[3873] =17;
weight[3874] =16;
weight[3875] =15;
weight[3876] =14;
weight[3877] =13;
weight[3878] =12;
weight[3879] =11;
weight[3880] =10;
weight[3881] =9;
weight[3882] =8;
weight[3883] =7;
weight[3884] =6;
weight[3885] =5;
weight[3886] =4;
weight[3887] =3;
weight[3888] =4;
weight[3889] =5;
weight[3890] =6;
weight[3891] =7;
weight[3892] =8;
weight[3893] =9;
weight[3894] =10;
weight[3895] =11;
weight[3896] =12;
weight[3897] =13;
weight[3898] =14;
weight[3899] =15;
weight[3900] =16;
weight[3901] =17;
weight[3902] =18;
weight[3903] =999;
weight[3904] =999;
weight[3905] =33;
weight[3906] =34;
weight[3907] =35;
weight[3908] =36;
weight[3909] =37;
weight[3910] =38;
weight[3911] =39;
weight[3912] =40;
weight[3913] =40;
weight[3914] =39;
weight[3915] =38;
weight[3916] =37;
weight[3917] =36;
weight[3918] =35;
weight[3919] =34;
weight[3920] =33;
weight[3921] =32;
weight[3922] =31;
weight[3923] =30;
weight[3924] =29;
weight[3925] =28;
weight[3926] =27;
weight[3927] =26;
weight[3928] =25;
weight[3929] =24;
weight[3930] =23;
weight[3931] =22;
weight[3932] =21;
weight[3933] =20;
weight[3934] =19;
weight[3935] =18;
weight[3936] =17;
weight[3937] =16;
weight[3938] =15;
weight[3939] =14;
weight[3940] =13;
weight[3941] =12;
weight[3942] =11;
weight[3943] =10;
weight[3944] =9;
weight[3945] =8;
weight[3946] =7;
weight[3947] =6;
weight[3948] =5;
weight[3949] =4;
weight[3950] =3;
weight[3951] =2;
weight[3952] =3;
weight[3953] =4;
weight[3954] =5;
weight[3955] =6;
weight[3956] =7;
weight[3957] =8;
weight[3958] =9;
weight[3959] =10;
weight[3960] =11;
weight[3961] =12;
weight[3962] =13;
weight[3963] =14;
weight[3964] =15;
weight[3965] =16;
weight[3966] =17;
weight[3967] =999;
weight[3968] =999;
weight[3969] =34;
weight[3970] =35;
weight[3971] =36;
weight[3972] =37;
weight[3973] =38;
weight[3974] =39;
weight[3975] =40;
weight[3976] =40;
weight[3977] =39;
weight[3978] =38;
weight[3979] =37;
weight[3980] =36;
weight[3981] =35;
weight[3982] =34;
weight[3983] =33;
weight[3984] =32;
weight[3985] =31;
weight[3986] =30;
weight[3987] =29;
weight[3988] =28;
weight[3989] =27;
weight[3990] =26;
weight[3991] =25;
weight[3992] =24;
weight[3993] =23;
weight[3994] =22;
weight[3995] =21;
weight[3996] =20;
weight[3997] =19;
weight[3998] =18;
weight[3999] =17;
weight[4000] =16;
weight[4001] =15;
weight[4002] =14;
weight[4003] =13;
weight[4004] =12;
weight[4005] =11;
weight[4006] =10;
weight[4007] =9;
weight[4008] =8;
weight[4009] =7;
weight[4010] =6;
weight[4011] =5;
weight[4012] =4;
weight[4013] =3;
weight[4014] =2;
weight[4015] =1;
weight[4016] =2;
weight[4017] =3;
weight[4018] =4;
weight[4019] =5;
weight[4020] =6;
weight[4021] =7;
weight[4022] =8;
weight[4023] =9;
weight[4024] =10;
weight[4025] =11;
weight[4026] =12;
weight[4027] =13;
weight[4028] =14;
weight[4029] =15;
weight[4030] =16;
weight[4031] =999;
weight[4032] =999;
weight[4033] =999;
weight[4034] =999;
weight[4035] =999;
weight[4036] =999;
weight[4037] =999;
weight[4038] =999;
weight[4039] =999;
weight[4040] =999;
weight[4041] =999;
weight[4042] =999;
weight[4043] =999;
weight[4044] =999;
weight[4045] =999;
weight[4046] =999;
weight[4047] =999;
weight[4048] =999;
weight[4049] =999;
weight[4050] =999;
weight[4051] =999;
weight[4052] =999;
weight[4053] =999;
weight[4054] =999;
weight[4055] =999;
weight[4056] =999;
weight[4057] =999;
weight[4058] =999;
weight[4059] =999;
weight[4060] =999;
weight[4061] =999;
weight[4062] =999;
weight[4063] =999;
weight[4064] =999;
weight[4065] =999;
weight[4066] =999;
weight[4067] =999;
weight[4068] =999;
weight[4069] =999;
weight[4070] =999;
weight[4071] =999;
weight[4072] =999;
weight[4073] =999;
weight[4074] =999;
weight[4075] =999;
weight[4076] =999;
weight[4077] =999;
weight[4078] =999;
weight[4079] =0;
weight[4080] =999;
weight[4081] =999;
weight[4082] =999;
weight[4083] =999;
weight[4084] =999;
weight[4085] =999;
weight[4086] =999;
weight[4087] =999;
weight[4088] =999;
weight[4089] =999;
weight[4090] =999;
weight[4091] =999;
weight[4092] =999;
weight[4093] =999;
weight[4094] =999;
weight[4095] =999;
end 
endmodule